* SPICE3 file created from SenseAmplifier.ext - technology: scmos

.include osu018.lib
.option scale=0.1u

M1000 d se blbar vdd1 pfet w=8 l=2
+  ad=60 pd=44 as=40 ps=26
M1001 a_n6_n18# se gnd gnd nfet w=8 l=2
+  ad=120 pd=78 as=40 ps=26
M1002 vdd1 d a_n6_18# vdd1 pfet w=4 l=2
+  ad=40 pd=36 as=60 ps=44
M1003 d a_n6_18# vdd1 vdd1 pfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 d a_n6_18# a_n6_n18# gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1005 a_n6_n18# d a_n6_18# gnd nfet w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1006 bl se a_n6_18# vdd1 pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
C0 d vdd1 0.55fF
C1 se bl 0.05fF
C2 a_n6_18# se 0.18fF
C3 d a_n6_n18# 0.16fF
C4 blbar vdd1 0.12fF
C5 d blbar 0.06fF
C6 vdd1 bl 0.12fF
C7 a_n6_18# vdd1 0.66fF
C8 a_n6_18# d 0.33fF
C9 a_n6_18# a_n6_n18# 0.16fF
C10 se vdd1 0.28fF
C11 d se 0.16fF
C12 se a_n6_n18# 0.20fF
C13 se blbar 0.05fF
C14 a_n6_18# bl 0.06fF
C15 a_n6_n18# gnd 0.12fF
C16 d gnd 0.25fF
C17 blbar gnd 0.00fF
C18 bl gnd 0.00fF
C19 a_n6_18# gnd 0.15fF
C20 se gnd 0.19fF
C21 vdd1 gnd 1.35fF
v3 vdd1 gnd  dc 1.8V
v2  bl gnd pulse(1.5V 1.5V 0ns 1ns 1ns 10ns 20ns)
v1  se gnd pulse(0V 1.8V 5ns 1ns 1ns 20ns 40ns)
v4  blbar gnd pulse(1.8V 1.8V 0ns 1ns 1ns 10ns 20ns)
.tran 5e-12 200e-09 0e-09

* Control Statements 
.control
run
plot bl blbar-2 se-4 d-6
.endc
.end
