* SPICE3 file created from Pre-Charge.ext - technology: scmos

.include osu018.lib
.option scale=0.1u

M1000 vdd2 pclk blbar w_n22_n11# pfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 blbar pclk bl w_n22_n11# pfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1002 vdd1 pclk bl w_n22_n11# pfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 pclk vdd1 0.05fF
C1 vdd2 w_n22_n11# 0.03fF
C2 pclk vdd2 0.05fF
C3 vdd2 blbar 0.04fF
C4 w_n22_n11# bl 0.09fF
C5 vdd1 bl 0.04fF
C6 w_n22_n11# vdd1 0.03fF
C7 pclk w_n22_n11# 0.34fF
C8 bl blbar 0.04fF
C9 w_n22_n11# blbar 0.09fF
v1 vdd1 gnd  dc 1.8V
v3 vdd2 gnd  dc 1.8V
v2  pclk gnd pulse(0 1.8V 0.1ns 1ns 1ns 30ns 60ns)
.tran 2e-12 100e-09 0e-09

* Control Statements 
.control
run
plot pclk bl-2 blbar-4
.endc
.end
